`include "../inc/defines.v"

module regfile (
        input   wire    rst,
        input   wire    clk,

        input   wire                    we,
        input   wire[`RegAddrBus]       waddr,
        input   wire[`RegBus]           wdata,

        input   wire                    re1,
        input   wire[`RegAddrBus]       raddr1,
        output  reg[`RegBus]            rdata1,

        input   wire                    re2,
        input   wire[`RegAddrBus]       raddr2,
        output  reg[`RegBus]            rdata2
);

reg[`RegBus]    regs[0:`RegNum-1];

// Write regisers
always @(posedge clk) begin
        if(rst == `RstDisable) begin
                if( (we == `WriteEnable) && (waddr != `RegNumLog2'h0) ) begin
                        regs[waddr] <= wdata;
                end
        end

end

// Read registers 1
always @(*) begin
        if(rst == `RstEnable) begin
                rdata1 = `ZeroWord;
        end else if(raddr1 == `RegNumLog2'h0) begin
                rdata1 = `ZeroWord;
        end else if( (raddr1 == waddr) && (we == `WriteEnable) && (re1 == `ReadEnable) ) begin
                // The 4th instruction want to read data from register x in decode stage,
                // but the data will write to the register in writeback stage(the next clk rising) by the first instruction.
                // So, we direct copy the write data to read data.
                rdata1 = wdata;
        end else if(re1 == `ReadEnable) begin
                rdata1 = regs[raddr1];
        end else begin
                rdata1 = `ZeroWord;
        end
end

// Read registers 2
always @(*) begin
        if(rst == `RstEnable) begin
                rdata2 = `ZeroWord;
        end else if(raddr2 == `RegNumLog2'h0) begin
                rdata2 = `ZeroWord;
        end else if( (raddr2 == waddr) && (we == `WriteEnable) && (re2 == `ReadEnable) ) begin
                // Same with 'read register 1'
                rdata2 = wdata;
        end else if(re2 == `ReadEnable) begin
                rdata2 = regs[raddr2];
        end else begin
                rdata2 = `ZeroWord;
        end
end


endmodule